// Copyright (c) 2024 Ethan Sifferman.
// All rights reserved. Distribution Prohibited.

// https://vesa.org/vesa-standards/
// http://tinyvga.com/vga-timing
module vga_timer (
    // TODO
    // possible ports list:
    // input  logic       clk_i,
    // input  logic       rst_ni,
    // output logic       hsync_o,
    // output logic       vsync_o,
    // output logic       visible_o,
    // output logic [8:0] position_x_o,
    // output logic [7:0] position_y_o
);

// TODO

endmodule
